module test_cpu_table32;
  top_node node_inst;

  initial begin
    node_inst  = new("top", null);
  end

endmodule
